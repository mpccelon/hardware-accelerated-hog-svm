module xillyvga_core
  (
  input  S_AXI_ACLK,
  input [31:0] S_AXI_ARADDR,
  input  S_AXI_ARESETN,
  input  S_AXI_ARVALID,
  input [31:0] S_AXI_AWADDR,
  input  S_AXI_AWVALID,
  input  S_AXI_BREADY,
  input  S_AXI_RREADY,
  input [31:0] S_AXI_WDATA,
  input [3:0] S_AXI_WSTRB,
  input  S_AXI_WVALID,
  input  clk_in,
  input  m_axi_aclk,
  input  m_axi_aresetn,
  input  m_axi_arready,
  input  m_axi_awready,
  input [1:0] m_axi_bresp,
  input  m_axi_bvalid,
  input [31:0] m_axi_rdata,
  input  m_axi_rlast,
  input [1:0] m_axi_rresp,
  input  m_axi_rvalid,
  input  m_axi_wready,
  output  S_AXI_ARREADY,
  output  S_AXI_AWREADY,
  output [1:0] S_AXI_BRESP,
  output  S_AXI_BVALID,
  output [31:0] S_AXI_RDATA,
  output [1:0] S_AXI_RRESP,
  output  S_AXI_RVALID,
  output  S_AXI_WREADY,
  output [31:0] m_axi_araddr,
  output [1:0] m_axi_arburst,
  output [3:0] m_axi_arcache,
  output [3:0] m_axi_arlen,
  output [2:0] m_axi_arprot,
  output [2:0] m_axi_arsize,
  output  m_axi_arvalid,
  output [31:0] m_axi_awaddr,
  output [1:0] m_axi_awburst,
  output [3:0] m_axi_awcache,
  output [3:0] m_axi_awlen,
  output [2:0] m_axi_awprot,
  output [2:0] m_axi_awsize,
  output  m_axi_awvalid,
  output  m_axi_bready,
  output  m_axi_rready,
  output [31:0] m_axi_wdata,
  output  m_axi_wlast,
  output [3:0] m_axi_wstrb,
  output  m_axi_wvalid,
  output vga_clk,
  output [7:0] vga_blue,
  output [7:0] vga_green,
  output  vga_hsync,
  output [7:0] vga_red,
  output  dvi_clk_n,
  output  dvi_clk_p,
  output [2:0] dvi_d_n,
  output [2:0] dvi_d_p,
  output  vga_de,
  output  vga_vsync
);
endmodule
